v1 4 0 10
vm 4 1 0
r1 1 2 2
r2 2 0 8
r3 2 3 4
f1 3 0 vm 3
i1 5 3 5
r4 5 0 6
r6 5 3 2

r1 a1 a 2
v1 a1 b 1
r3 c  d 4
t1 c d a b 10

r1 a a1 2
v1 a 0 1
r3 c  0 4
t1 a1 0 c 0 10

vsrc1 a 0 0
f2 e 0 vsrc1 2 
isrc3 a 0 4
r4  e 0 5

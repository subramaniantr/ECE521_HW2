vsrc2 a 0 5
e1 c 0 a 0 2
r3 c 0 10

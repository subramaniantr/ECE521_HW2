r1 a1 a 2
v1 a1 0 1
r3 c  0 4
Nt1 a 0 c 0 10

v1 4 0 24
vm 4 1 0
r1 1 2 10
r2 2 0 12
r3 4 3 24
r4 2 3 4
h1 3 0 vm 4

v1 a 0 1
r3 c  0 4
t1 c 0 a 0 10

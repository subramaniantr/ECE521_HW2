v1 a b 1
r3 c 0 4
Ot1 c a b 10

r2 node4 1 100
r3 1 2 100
r4 2 3 100
r5 3 0 100
v1 node4 0 10

vsrc2 a b 5
e1 c d a b 2
r3 c d 10

v1 c 0 5
g3 a 0 c 0 3 
r1 a 0 10

g3 h i j k 3 

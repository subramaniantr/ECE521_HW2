r1      1                                3                           1.0
d1 1 2    dmod 2.0


d3 2 3  dmod2 1
v2 3 0 5
d4 1 3  dmod 3
cyy 4 0 1e-12
v100 3 4 2.5
dfoo 3 2 dmod 1

m1 1 2 3 4 mmod 1          1
m2 2 3          3 0 mmod2 10 2
cxx 3 0 1e-12
mdiode          2 2 3 0 mmod 10 10

v1 1 0 1

r2 2 0 3.0
g1 1 2 3          4 2.0
r3 3      4 5.0

i1 2 0 3
i2 1 3 2.5

c1 2 3          3e-12


e1 1 2 3 4          1
h1          3 4 1 2 1.5
f1 3          4 2 0 5.5

v1 1 2 20
r1 1 0 2
r2 2 3 6
r3 3 0 4
r4 1 4 3
r5 4 0 1
i1 0 2 10
e1 3 4 1 4 3

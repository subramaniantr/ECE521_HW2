vsrc1 a b 0
h4 c d vsrc1 4 
isrc3 a b 2
r4  c d 5

v1 a 0 1
r3 c 0 4
Ot1 a 0 c 10
